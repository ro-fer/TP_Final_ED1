-- Contador de unos

-- Estudiante: Fernandez, Rocio

library IEEE;
use IEEE.std_logic_1164.all;
